library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top_level_tb is
end;

architecture a_top_level_tb of top_level_tb is
    component fetch is port (
        clk                 : in std_logic;
        rst                 : in std_logic;
        pc_wr_en            : in std_logic;
        rd_rom              : in std_logic;
        instruction         : out unsigned(15 downto 0)
    );
    end component;

    component decode is port (
        clk             : in std_logic;
        rst             : in std_logic;
        instruction     : in unsigned(15 downto 0);
        rd_rom          : out std_logic;
        operation       : out unsigned(1 downto 0)
    );
    end component;

    component execute is port (
        clk             : in std_logic;
        rst             : in std_logic;
        entr0           : in unsigned(15 downto 0);
        entr1           : in unsigned(15 downto 0);
        operation       : in unsigned(1 downto 0);
        result          : out unsigned(15 downto 0)
    );
    end component;

    constant period_time            : time := 100 ns;
    signal finished                 : std_logic := '0';
    signal clk, rst                 : std_logic;
    signal pc_wr_en, rd_rom         : std_logic;
    signal instruction, result      : unsigned(15 downto 0);
    signal operation                : unsigned(1 downto 0);

begin

    fetch_uut : fetch port map(
        clk => clk,
        rst => rst,
        pc_wr_en => pc_wr_en,
        rd_rom => rd_rom,
        instruction => instruction
    );

    decode_uut : decode port map(
        clk => clk,
        rst => rst,
        rd_rom => rd_rom,
        instruction => instruction,
        operation => operation
    );

    execute_uut : execute port map(
        clk => clk,
        rst => rst,
        entr0 => instruction,
        entr1 => instruction,
        operation => operation,
        result => result
    );

    reset_global: process
    begin
        rst <= '1';
        wait for period_time*2;
        rst <= '0';
        wait;
    end process;

    sim_time_proc: process
    begin
        wait for 10 us;         -- <== TEMPO TOTAL DA SIMULACAO!!!
        finished <= '1';
        wait;
    end process sim_time_proc;

    clk_proc: process
    begin                       -- gera clock até que sim_time_proc termine
        while finished /= '1' loop
            clk <= '0';
            wait for period_time/2;
            clk <= '1';
            wait for period_time/2;
        end loop;
        wait;
    end process clk_proc;

    process
    begin
        wait for 200 ns;
        pc_wr_en <= '1';

        wait;
    end process;
end architecture;