library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fetch_tb is
end;

architecture a_fetch_tb of fetch_tb is
    component fetch is port (
        clk                 : in std_logic;
        rst                 : in std_logic;
        pc_wr_en            : in std_logic
    );
    end component;

    constant period_time            : time := 100 ns;
    signal finished                 : std_logic := '0';
    signal clk, rst                 : std_logic;
    signal pc_wr_en      : std_logic;

begin

    fetch_uut : fetch port map(
        clk => clk,
        rst => rst,
        pc_wr_en => pc_wr_en
    );

    reset_global: process
    begin
        rst <= '1';
        wait for period_time*2;
        rst <= '0';
        wait;
    end process;

    sim_time_proc: process
    begin
        wait for 10 us;         -- <== TEMPO TOTAL DA SIMULACAO!!!
        finished <= '1';
        wait;
    end process sim_time_proc;

    clk_proc: process
    begin                       -- gera clock até que sim_time_proc termine
        while finished /= '1' loop
            clk <= '0';
            wait for period_time/2;
            clk <= '1';
            wait for period_time/2;
        end loop;
        wait;
    end process clk_proc;

    process
    begin
        wait for 200 ns;
        pc_wr_en <= '1';

        wait;
    end process;
end architecture;