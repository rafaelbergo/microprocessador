library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port (
        clk:        in std_logic;
        address:    in unsigned(6 downto 0);
        data:       out unsigned(16 downto 0);
        rd_rom:     in std_logic
    );
end entity;

-- OPCODES:

-- 0000 NOP
-- 0001 SW
-- 0010 LD
-- 0011 MOV (A,R) or (R,A)
-- 0100 ADD
-- 0101 SUBI
-- 0110 SUB
-- 0111 LW
-- 1000 MOV (R,R)
-- 1001 BLE
-- 1010 JUMP
-- 1011 BLO
-- 1100 CMPR
-- 1101 AND
-- 1110 OR
-- 1111

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(16 downto 0);
    constant content_rom: mem := (
         -- INICIALIZACAO
        0   =>  B"0010_0_0000_00000010", -- LD R0,2
        1   =>  B"0010_0_0001_00000001", -- LD R1,1
        2   =>  B"0010_0_0011_00000010", -- LD R3,2
        3   =>  B"0010_0_0100_00000100", -- LD R4,4
        4   =>  B"0010_0_1000_00000000", -- LD R8,0
        5   =>  B"0011_1_0000_00000000", -- MOV A,R0

         -- POPULA OS 32 PRIMEIROS BITS
        6   =>  B"0001_0_0000_00000000", -- SW A,0(R0)
        7   =>  B"0100_0_0001_00000000", -- ADD A,R1
        8   =>  B"0011_0_0000_00000000", -- MOV R0,A
        9   =>  B"0101_0_0000_00100000", -- SUBI A,32
        10  =>  B"1001_0_0000_11111010", -- BLE -5
        11  =>  B"1010_0_0000_00010011", -- JUMP 19

         -- ZERA O NUMERO NAO PRIMO
        12  =>  B"0011_1_1000_00000000", -- MOV A,R8
        13  =>  B"0001_0_0100_00000000", -- SW A,0(R4)
        14  =>  B"1010_0_0000_00011000", -- JUMP 24

         -- FUNCAO QUE DIVIDE
        15  =>  B"0110_0_0101_00000000", -- SUB A,R5
        16  =>  B"1011_0_0000_00000111", -- BLO 7
        17  =>  B"1001_0_0000_11111010", -- BLE -6
        18  =>  B"1010_0_0000_00001111", -- JUMP 15

        -- LOOP PRINCIPAL
        19  =>  B"0111_0_0011_00000000", -- LW A,0(R3)
        20  =>  B"0001_0_1000_00100011", -- SW A,35(R8)
        21  =>  B"0011_0_0101_00000000", -- MOV R5,A
        22  =>  B"0111_0_0100_00000000", -- LW A,0(R4)
        23  =>  B"1010_0_0000_00001111", -- JUMP 15 (FUNCAO DIVISAO)

        -- INCREMENTA R4
        24  =>  B"0011_1_0100_00000000", -- MOV A,R4
        25  =>  B"0100_0_0001_00000000", -- ADD A,R1
        26  =>  B"0011_0_0100_00000000", -- MOV R4,A
        27  =>  B"0101_0_0000_00100000", -- SUBI A,32
        28  =>  B"1001_0_0000_11111001", -- BLE -7

        -- INCREMETA R3
        29  =>  B"0011_1_0011_00000000", -- MOV A,R3
        30  =>  B"0100_0_0001_00000000", -- ADD A,R1
        31  =>  B"0011_0_0011_00000000", -- MOV R3,A
        32  =>  B"0101_0_0000_00100000", -- SUBI A,32
        33  =>  B"1011_0_0000_00000001", -- BLO 1
        34  =>  B"1010_0_0000_00101011", -- JUMP 43 (SAI DO LOOP)
        35  =>  B"0111_0_0011_00000000", -- LW A,0(R3)
        36  =>  B"0101_0_0000_00000000", -- SUBI A,0 (VERIFICA SE O CONTEUDO NAO E 0)
        37  =>  B"1001_0_0000_11110111", -- BLE -9
        38  =>  B"0011_1_0011_00000000", -- MOV A,R3
        39  =>  B"0100_0_0001_00000000", -- ADD A,R1
        40  =>  B"0100_0_0001_00000000", -- ADD A,R1
        41  =>  B"0011_0_0100_00000000", -- MOV R4,A
        42  =>  B"1010_0_0000_00010011", -- JUMP 19

        -- CARREGA 1171 NO ACUMULADOR
        43  =>  B"0011_1_1000_00000000", -- MOV A,R8
        44  =>  B"0001_0_1000_00100100", -- SW A,36(R8)
        45  =>  B"0010_0_0000_01111111", -- LD R0,127
        46  =>  B"0011_1_0000_00000000", -- MOV A,R0
        47  =>  B"0100_0_0000_00000000", -- ADD A,R0
        48  =>  B"0011_0_0000_00000000", -- MOV R0,A
        49  =>  B"0100_0_0000_00000000", -- ADD A,R0
        50  =>  B"0011_0_0000_00000000", -- MOV R0,A
        51  =>  B"0100_0_0000_00000000", -- ADD A,R0
        52  =>  B"0010_0_0000_01111111", -- LD R0,127
        53  =>  B"0100_0_0000_00000000", -- ADD A,R0
        54  =>  B"0010_0_0000_00011100", -- LD R0,28
        55  =>  B"0100_0_0000_00000000", -- ADD A,R0
        56  =>  B"0001_0_0100_00000000", -- SW A,0(R4)
        57  =>  B"0010_0_0011_00000010", -- LD R3,2
        58  =>  B"1010_0_0000_01000001", -- JUMP 65

        59  =>  B"0011_1_0011_00000000", -- MOV A,R3
        60  =>  B"0100_0_0001_00000000", -- ADD A,R1
        61  =>  B"0011_0_0011_00000000", -- MOV R3,A
        62  =>  B"0101_0_0000_00100000", -- SUBI A,32
        63  =>  B"1001_0_0000_00000001", -- BLE 1
        64  =>  B"1010_0_0000_01001010", -- JUMP 74
        
        65  =>  B"0111_0_0011_00000000", -- LW A,0(R3)
        66  =>  B"0101_0_0000_00000000", -- SUBI A,0
        67  =>  B"1001_0_0000_11110111", -- BLE -9
        68  =>  B"0011_0_0101_00000000", -- MOV R5,A
        69  =>  B"0111_0_0100_00000000", -- LW A,0(R4)

        70  =>  B"0110_0_0101_00000000", -- SUB A,R5
        71  =>  B"1011_0_0000_11110011", -- BLO -13
        72  =>  B"1001_0_0000_00000011", -- BLE 3
        73  =>  B"1010_0_0000_01000110", -- JUMP 70
        
        74  =>  B"0011_1_0001_00000000", -- MOV A,R1
        75  =>  B"0001_0_1000_00100100", -- SW A,36(R8)
        others => (others => '0')
    );
begin
    process(clk)
    begin
        if rising_edge(clk) and rd_rom = '1' then 
            data <= content_rom(to_integer(address));
        end if;
    end process;
end architecture;